library ieee ;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

entity Pong is
  port (
    MAX10_CLK1_50 : in std_logic;
    
  ) ;
end Pong ;

architecture work of Pong is



begin



end architecture ; -- work